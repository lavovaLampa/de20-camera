package vga_pkg is
    constant IMG_HEIGHT : natural := 480;
    constant IMG_WIDTH  : natural := 640;

    constant HBLANK_PIXELS : natural := 160;
    constant VBLANK_LINES  : natural := 44;
end package vga_pkg;
