library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity project_top is
    port(
        clk : in std_logic;
        rst : in std_logic
    );
end entity project_top;

architecture RTL of project_top is
    
begin

end architecture RTL;
